module JKFF(output Q,q,input J,K,clk);//jkflip-flop

wire x,y,Q,q;




and a1(x,K,Q,clk);
and a2(y,J,q,clk);
nor n1(Q,q,x);
nor n2(q,Q,y);
endmodule
